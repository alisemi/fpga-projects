`timescale 1ns / 1ps

module MatrixDriver(
    input logic clk,
    input logic [5:0] letter,
    output logic oe, //output enable	
    output logic SH_CP, // shift register clk pulse
    output logic ST_CP, // store register clk pulse
    output logic reset, // reset for the shift register
    output logic DS, // digital signal
    output logic [7:0] row);
        
    // message ve row buradan matrix modulune verilecek
    logic [7:0][23:0] data;
    
    always_ff@(posedge clk)
        case(letter)
            6'b000_000: begin // D_START
                data[0] <= 24'b00000000_00000000_11111111;
                data[1] <= 24'b00000000_00000000_11111111;
                data[2] <= 24'b00000000_00000000_11111111;
                data[3] <= 24'b00000000_00000000_11111111;
                data[4] <= 24'b00000000_00000000_11111111;
                data[5] <= 24'b00000000_00000000_11111111;
                data[6] <= 24'b00000000_00000000_11111111;
                data[7] <= 24'b00000000_00000000_11111111;
            end
            6'b000_001: begin // A
                data[0] <= 24'b00111100_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11111111_00000000_00000000;
                data[6] <= 24'b11000011_00000000_00000000;
                data[7] <= 24'b11000011_00000000_00000000;
            end
            6'b000_010: begin // B
                data[0] <= 24'b11111110_00000000_00000000;
                data[1] <= 24'b11000001_00000000_00000000;
                data[2] <= 24'b11000001_00000000_00000000;
                data[3] <= 24'b11111110_00000000_00000000;
                data[4] <= 24'b11111110_00000000_00000000;
                data[5] <= 24'b11000001_00000000_00000000;
                data[6] <= 24'b11000001_00000000_00000000;
                data[7] <= 24'b11111110_00000000_00000000;
            end
            6'b000_011: begin // C
                data[0] <= 24'b01111100_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000000_00000000_00000000;
                data[4] <= 24'b11000000_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b01111100_00000000_00000000;
            end
            6'b000_100: begin // D
                data[0] <= 24'b11111100_00000000_00000000;
                data[1] <= 24'b11111110_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11000011_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b11111110_00000000_00000000;
                data[7] <= 24'b01111100_00000000_00000000;
            end
            6'b000_101: begin // E
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11111111_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11000000_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b000_110: begin // F
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11111000_00000000_00000000;
                data[4] <= 24'b11111000_00000000_00000000;
                data[5] <= 24'b11000000_00000000_00000000;
                data[6] <= 24'b11000000_00000000_00000000;
                data[7] <= 24'b11000000_00000000_00000000;
            end
            6'b000_111: begin // G
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11011111_00000000_00000000;
                data[4] <= 24'b11011111_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b001_000: begin // H
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11000011_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11111111_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b11000011_00000000_00000000;
                data[7] <= 24'b11000011_00000000_00000000;
            end
            6'b001_001: begin // I
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b00011000_00000000_00000000;
                data[3] <= 24'b00011000_00000000_00000000;
                data[4] <= 24'b00011000_00000000_00000000;
                data[5] <= 24'b00011000_00000000_00000000;
                data[6] <= 24'b01111110_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b001_010: begin // J
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b00011000_00000000_00000000;
                data[3] <= 24'b00011000_00000000_00000000;
                data[4] <= 24'b00011000_00000000_00000000;
                data[5] <= 24'b00011000_00000000_00000000;
                data[6] <= 24'b01111000_00000000_00000000;
                data[7] <= 24'b01111000_00000000_00000000;
            end
            6'b001_011: begin // K
                data[0] <= 24'b0011_0001_0000000000000000;
                data[1] <= 24'b0011_0011_0000000000000000;
                data[2] <= 24'b0011_0110_0000000000000000;
                data[3] <= 24'b0011_1100_0000000000000000;
                data[4] <= 24'b0011_1100_0000000000000000;
                data[5] <= 24'b0011_0110_0000000000000000;
                data[6] <= 24'b0011_0011_0000000000000000;
                data[7] <= 24'b0011_0001_0000000000000000;
            end
            6'b001_100: begin // L
                data[0] <= 24'b11000000_00000000_00000000;
                data[1] <= 24'b11000000_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11000000_00000000_00000000;
                data[4] <= 24'b11000000_00000000_00000000;
                data[5] <= 24'b11000000_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b001_101: begin // M
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11100111_00000000_00000000;
                data[2] <= 24'b11111111_00000000_00000000;
                data[3] <= 24'b10011001_00000000_00000000;
                data[4] <= 24'b10000001_00000000_00000000;
                data[5] <= 24'b10000001_00000000_00000000;
                data[6] <= 24'b10000001_00000000_00000000;
                data[7] <= 24'b10000001_00000000_00000000;
            end
            6'b001_110: begin // N
                data[0] <= 24'b11000001_00000000_00000000;
                data[1] <= 24'b11100001_00000000_00000000;
                data[2] <= 24'b10110001_00000000_00000000;
                data[3] <= 24'b10011001_00000000_00000000;
                data[4] <= 24'b10001101_00000000_00000000;
                data[5] <= 24'b10000111_00000000_00000000;
                data[6] <= 24'b10000011_00000000_00000000;
                data[7] <= 24'b10000001_00000000_00000000;
            end
            6'b001_111: begin // O
                data[0] <= 24'b00111100_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11000011_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b01111110_00000000_00000000;
                data[7] <= 24'b00111100_00000000_00000000;
            end
            6'b010_000: begin // P
                data[0] <= 24'b11111000_00000000_00000000;
                data[1] <= 24'b11111100_00000000_00000000;
                data[2] <= 24'b11000110_00000000_00000000;
                data[3] <= 24'b11000110_00000000_00000000;
                data[4] <= 24'b11111100_00000000_00000000;
                data[5] <= 24'b11111000_00000000_00000000;
                data[6] <= 24'b11000000_00000000_00000000;
                data[7] <= 24'b11000000_00000000_00000000;
            end
            6'b010_001: begin // Q
                data[0] <= 24'b00111100_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11000011_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b01111100_00000000_00000000;
                data[7] <= 24'b00111111_00000000_00000000;
            end
            6'b010_010: begin // R
                data[0] <= 24'b11111000_00000000_00000000;
                data[1] <= 24'b10001100_00000000_00000000;
                data[2] <= 24'b10001100_00000000_00000000;
                data[3] <= 24'b10001100_00000000_00000000;
                data[4] <= 24'b11111000_00000000_00000000;
                data[5] <= 24'b10001000_00000000_00000000;
                data[6] <= 24'b10000100_00000000_00000000;
                data[7] <= 24'b10000010_00000000_00000000;
            end
            6'b010_011: begin // S
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11111110_00000000_00000000;
                data[4] <= 24'b01111111_00000000_00000000;
                data[5] <= 24'b00000011_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b010_100: begin // T
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b00011000_00000000_00000000;
                data[3] <= 24'b00011000_00000000_00000000;
                data[4] <= 24'b00011000_00000000_00000000;
                data[5] <= 24'b00011000_00000000_00000000;
                data[6] <= 24'b00011000_00000000_00000000;
                data[7] <= 24'b00011000_00000000_00000000;
            end
            6'b010_101: begin // U
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11000011_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11000011_00000000_00000000;
                data[5] <= 24'b11000011_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b010_110: begin // V
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11000011_00000000_00000000;
                data[2] <= 24'b11000011_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11000011_00000000_00000000;
                data[5] <= 24'b01111110_00000000_00000000;
                data[6] <= 24'b00111100_00000000_00000000;
                data[7] <= 24'b00011000_00000000_00000000;
            end
            6'b010_111: begin // W
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11000011_00000000_00000000;
                data[2] <= 24'b11011011_00000000_00000000;
                data[3] <= 24'b11011011_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11100111_00000000_00000000;
                data[6] <= 24'b11000011_00000000_00000000;
                data[7] <= 24'b11000011_00000000_00000000;
            end
            6'b011_000: begin // X
                data[0] <= 24'b11000011_00000000_00000000;
                data[1] <= 24'b11100111_00000000_00000000;
                data[2] <= 24'b01111110_00000000_00000000;
                data[3] <= 24'b00111100_00000000_00000000;
                data[4] <= 24'b00111100_00000000_00000000;
                data[5] <= 24'b01111110_00000000_00000000;
                data[6] <= 24'b11100111_00000000_00000000;
                data[7] <= 24'b11000011_00000000_00000000;
            end
            6'b011_001: begin // Y
                data[0] <= 24'b11100111_00000000_00000000;
                data[1] <= 24'b11100111_00000000_00000000;
                data[2] <= 24'b11100111_00000000_00000000;
                data[3] <= 24'b11100111_00000000_00000000;
                data[4] <= 24'b00111100_00000000_00000000;
                data[5] <= 24'b00111100_00000000_00000000;
                data[6] <= 24'b00111100_00000000_00000000;
                data[7] <= 24'b00111100_00000000_00000000;
            end
            6'b011_010: begin // Z
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b00001110_00000000_00000000;
                data[3] <= 24'b00011100_00000000_00000000;
                data[4] <= 24'b00111000_00000000_00000000;
                data[5] <= 24'b01110000_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b100_000: begin // D0
                data[0] <= 24'b00111100_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b01100110_00000000_00000000;
                data[3] <= 24'b01100110_00000000_00000000;
                data[4] <= 24'b01100110_00000000_00000000;
                data[5] <= 24'b01100110_00000000_00000000;
                data[6] <= 24'b01111110_00000000_00000000;
                data[7] <= 24'b00111100_00000000_00000000;
            end
            6'b100_001: begin // D1
                data[0] <= 24'b00111000_00000000_00000000;
                data[1] <= 24'b01111000_00000000_00000000;
                data[2] <= 24'b01011000_00000000_00000000;
                data[3] <= 24'b00011000_00000000_00000000;
                data[4] <= 24'b00011000_00000000_00000000;
                data[5] <= 24'b00011000_00000000_00000000;
                data[6] <= 24'b01111110_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b100_010: begin // D2
                data[0] <= 24'b00111100_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000111_00000000_00000000;
                data[3] <= 24'b00001110_00000000_00000000;
                data[4] <= 24'b00011100_00000000_00000000;
                data[5] <= 24'b00111000_00000000_00000000;
                data[6] <= 24'b01110000_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b100_011: begin // D3
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b01111110_00000000_00000000;
                data[2] <= 24'b00000110_00000000_00000000;
                data[3] <= 24'b00011110_00000000_00000000;
                data[4] <= 24'b00011110_00000000_00000000;
                data[5] <= 24'b00000110_00000000_00000000;
                data[6] <= 24'b01111110_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b100_100: begin // D4
                data[0] <= 24'b11000000_00000000_00000000;
                data[1] <= 24'b11000000_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11000011_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11111111_00000000_00000000;
                data[6] <= 24'b00000011_00000000_00000000;
                data[7] <= 24'b00000011_00000000_00000000;
            end
            6'b100_101: begin // D5
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11000000_00000000_00000000;
                data[3] <= 24'b11111111_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b00000011_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            6'b100_110: begin // D6
                data[0] <= 24'b01111000_00000000_00000000;
                data[1] <= 24'b01111000_00000000_00000000;
                data[2] <= 24'b01100000_00000000_00000000;
                data[3] <= 24'b01100000_00000000_00000000;
                data[4] <= 24'b01111110_00000000_00000000;
                data[5] <= 24'b01100110_00000000_00000000;
                data[6] <= 24'b01100110_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b100_111: begin // D7
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b00000110_00000000_00000000;
                data[3] <= 24'b00001100_00000000_00000000;
                data[4] <= 24'b00011000_00000000_00000000;
                data[5] <= 24'b00110000_00000000_00000000;
                data[6] <= 24'b01100000_00000000_00000000;
                data[7] <= 24'b11000000_00000000_00000000;
            end
            6'b101_000: begin // D8
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b01000010_00000000_00000000;
                data[2] <= 24'b01111110_00000000_00000000;
                data[3] <= 24'b00111100_00000000_00000000;
                data[4] <= 24'b00111100_00000000_00000000;
                data[5] <= 24'b01111110_00000000_00000000;
                data[6] <= 24'b01000010_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b101_001: begin // D9
                data[0] <= 24'b01111110_00000000_00000000;
                data[1] <= 24'b01000010_00000000_00000000;
                data[2] <= 24'b01000010_00000000_00000000;
                data[3] <= 24'b01000010_00000000_00000000;
                data[4] <= 24'b01111110_00000000_00000000;
                data[5] <= 24'b00000010_00000000_00000000;
                data[6] <= 24'b00000010_00000000_00000000;
                data[7] <= 24'b01111110_00000000_00000000;
            end
            6'b111_111: begin // INVALID
                data[0] <= 24'b00000000_11111111_00000000;
                data[1] <= 24'b00000000_11111111_00000000;
                data[2] <= 24'b00000000_11111111_00000000;
                data[3] <= 24'b00000000_11111111_00000000;
                data[4] <= 24'b00000000_11111111_00000000;
                data[5] <= 24'b00000000_11111111_00000000;
                data[6] <= 24'b00000000_11111111_00000000;
                data[7] <= 24'b00000000_11111111_00000000;
            end
            default: begin // Default
                data[0] <= 24'b11111111_00000000_00000000;
                data[1] <= 24'b11111111_00000000_00000000;
                data[2] <= 24'b11111111_00000000_00000000;
                data[3] <= 24'b11111111_00000000_00000000;
                data[4] <= 24'b11111111_00000000_00000000;
                data[5] <= 24'b11111111_00000000_00000000;
                data[6] <= 24'b11111111_00000000_00000000;
                data[7] <= 24'b11111111_00000000_00000000;
            end
            endcase
         
    DotMatrix dm(clk, data, oe, SH_CP, ST_CP, reset, DS, row);
        
endmodule
